library	IEEE;
use IEEE.STD_LOGIC_1164.all; 

package vectorul8 is
	type tip_matrice8 is array(15 downto 0) of std_logic_vector(7 downto 0);	
end package;  