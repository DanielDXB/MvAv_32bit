library	IEEE;
use IEEE.STD_LOGIC_1164.all; 

package vectorul4 is
	type tip_matrice4 is array(15 downto 0) of std_logic_vector(3 downto 0);	
end package;  